package shared_pkg;
    localparam MEM_DEPTH = 256;
    localparam ADDR_SIZE = $clog2(MEM_DEPTH);
endpackage